/* Copyright 2018 Tymoteusz Blazejczyk
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

/* Package: logic_unit_test_pkg
 *
 * Logic unit test package.
 */
package logic_unit_test_pkg;
`include "logic_avalon_st_driver_rx.svh"
`include "logic_avalon_st_driver_tx.svh"
`include "logic_axi4_stream_driver_rx.svh"
`include "logic_axi4_stream_driver_tx.svh"
`include "logic_axi4_lite_driver_slave.svh"
`include "logic_axi4_lite_driver_master.svh"
endpackage
