/* Copyright 2017 Tymoteusz Blazejczyk
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * @copyright
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

`ifndef LOGIC_AXI4_STREAM_SVH
`define LOGIC_AXI4_STREAM_SVH

`ifndef LOGIC_AXI4_STREAM_TDATA_BYTES
    `define LOGIC_AXI4_STREAM_TDATA_BYTES 1
`endif

`ifndef LOGIC_AXI4_STREAM_TID_WIDTH
    `define LOGIC_AXI4_STREAM_TID_WIDTH 1
`endif

`ifndef LOGIC_AXI4_STREAM_TDEST_WIDTH
    `define LOGIC_AXI4_STREAM_TDEST_WIDTH 1
`endif

`ifndef LOGIC_AXI4_STREAM_TUSER_WIDTH
    `define LOGIC_AXI4_STREAM_TUSER_WIDTH 1
`endif

`endif /* LOGIC_AXI4_STREAM_SVH */
