/* Copyright 2018 Tymoteusz Blazejczyk
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 */

`include "logic.svh"

/* Module: logic_axi4_stream_demux
 *
 * It will extract AXI4-Stream packets based on their unique tdest or tid
 * value from rx input to the second tx output. Remaning packets will be pass
 * through the first tx input.
 *
 * Parameters:
 *  PACKETS     - Number of packets with unique tdest (or tid) to extract
 *                from rx input to second tx output.
 *  EXTRACT     - List of unique packet identifiers tdest or tid.
 *  TDATA_BYTES - Number of bytes for tdata signal.
 *  TDEST_WIDTH - Number of bits for tdest signal.
 *  TUSER_WIDTH - Number of bits for tuser signal.
 *  TID_WIDTH   - Number of bits for tid signal.
 *  USE_TKEEP   - Enable or disable tkeep signal.
 *  USE_TSTRB   - Enable or disable tstrb signal.
 *  USE_TLAST   - Enable or disable tlast signal.
 *  USE_TID     - Use tid instead of tdest signal for extracting.
 *
 * Ports:
 *  aclk        - Clock.
 *  areset_n    - Asynchronous active-low reset.
 *  rx          - AXI4-Stream Rx interface.
 *  tx          - AXI4-Stream Tx interface. The second output is used for
 *                extracting packets from rx input based on EXTRACT list.
 */
module logic_axi4_stream_extract #(
    int PACKETS = 1,
    int TDATA_BYTES = 1,
    int TDEST_WIDTH = 1,
    int TUSER_WIDTH = 1,
    int TID_WIDTH = 1,
    int USE_TLAST = 1,
    int USE_TKEEP = 1,
    int USE_TSTRB = 1,
    int USE_TID = 1,
    int EXTRACT_WIDTH = (USE_TID > 0) ? TID_WIDTH : TUSER_WIDTH,
    bit [PACKETS-1:0][EXTRACT_WIDTH-1:0] EXTRACT = init_extract()
) (
    input aclk,
    input areset_n,
    `LOGIC_MODPORT(logic_axi4_stream_if, rx) rx,
    `LOGIC_MODPORT(logic_axi4_stream_if, tx) tx[2]
);
    typedef bit [PACKETS-1:0][EXTRACT_WIDTH-1:0] extract_t;

    function extract_t init_extract;
        for (int i = 0; i < PACKETS; ++i) begin
            init_extract[i] = i[EXTRACT_WIDTH-1:0];
        end
    endfunction

    logic areset_n_synced;

    logic_reset_synchronizer
    reset_synchronizer (
        .*
    );

    logic_axi4_stream_extract_main #(
        .PACKETS(PACKETS),
        .EXTRACT(EXTRACT),
        .TDATA_BYTES(TDATA_BYTES),
        .TDEST_WIDTH(TDEST_WIDTH),
        .TUSER_WIDTH(TUSER_WIDTH),
        .TID_WIDTH(TID_WIDTH),
        .USE_TLAST(USE_TLAST),
        .USE_TKEEP(USE_TKEEP),
        .USE_TSTRB(USE_TSTRB),
        .USE_TID(USE_TID)
    )
    main (
        .areset_n(areset_n_synced),
        .*
    );
endmodule
